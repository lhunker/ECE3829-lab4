`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:58:15 10/09/2014 
// Design Name: 
// Module Name:    lab4 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lab4(
    input [2:0] sw,
    input clk,
    input reset,
    output [6:0] seg,
    output [3:0] anode,
    output HS,
    output VS,
    output [2:0] red,
    output [2:0] grn,
    output [1:0] blu
    );


endmodule
